
module processor(
	input clock,
	input reset
);




